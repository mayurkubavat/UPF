module or_gate(output z, input x, y);

   assign z = x | y;

endmodule
